library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity sin_table is
port (
  i_clk          : in  std_logic;
  i_addr         : in  std_logic_vector(7 downto 0);
  o_data         : out std_logic_vector(11 downto 0));
end sin_table;
architecture rtl of sin_table is
type t_sin_table is array(0 to 199) of integer range -2048 to 2047;--range 0 to 4095;
constant C_SIN_TABLE  : t_sin_table := (
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633,
		 0,
	  633,
	 1204,
	 1657,
	 1948,
	 2047,
	 1948,
	 1657,
	 1204,
	  633,
		 0,
	 -633,
	-1204,
	-1657,
	-1948,
	-2048,
	-1948,
	-1657,
	-1204,
	 -633

--     2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415,
-- 2048,
-- 2681,
-- 3252,
-- 3705,
-- 3996,
-- 4095,
-- 3996,
-- 3705,
-- 3252,
-- 2681,
-- 2048,
-- 1415,
--  844,
--  391,
--  100,
--    0,
--  100,
--  391,
--  844,
-- 1415
);
begin
--------------------------------------------------------------------
p_table : process(i_clk)
begin
  if(rising_edge(i_clk)) then
    o_data  <= std_logic_vector(to_signed(C_SIN_TABLE(to_integer(unsigned(i_addr))),12));
  end if;
end process p_table;
end rtl;