library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;
use STD.textio.all;
use ieee.std_logic_textio.all;

library work;
use work.constants.all;
use work.records.all;
 
ENTITY Goertzel_tb IS
END Goertzel_tb;

ARCHITECTURE behavior OF Goertzel_tb IS 
	-- Component Declaration for the Unit Under Test (UUT)
	COMPONENT Goertzel is
	Port ( 	i_CLK : in  STD_LOGIC; -- Clock input
				i_ENABLE : in  STD_LOGIC; -- Enable input
				i_SIG : in  SIGNED(INPUT_WIDTH-1 downto 0); -- Signal 1
				i_COEFF : in SIGNED(CALC_WIDTH-1 downto 0); -- Coefficient input
				o_DFT : out  goertzel_result_type; -- DFT output
				o_NEW_RESULT : out  STD_LOGIC -- New result flag
			 );
	end COMPONENT;
	
	-- File
	file file_VECTORS : text;
	file file_RESULTS : text;
	constant c_WIDTH : natural := 4;
	constant signal_period : time := 2 us;
	-- Inputs
	signal i_CLK :  STD_LOGIC := '0'; -- Clock input
	signal i_ENABLE :  STD_LOGIC := '0'; -- Enable input
	signal i_SIG :  SIGNED(INPUT_WIDTH-1 downto 0) := (others => '0'); -- Signal 1
	signal i_COEFF : SIGNED(CALC_WIDTH-1 downto 0) := (others => '0'); -- Coefficient input
	-- Outputs
	signal o_DFT :  goertzel_result_type; -- DFT output
	signal o_NEW_RESULT : STD_LOGIC; -- New result flag
	
	-- Clock period definitions
   constant c_clk_period : time := 100 ns;

BEGIN
	-- Instantiate the Unit Under Test (UUT)
	uut: Goertzel PORT MAP( 	
				i_CLK => i_CLK,
				i_ENABLE => i_ENABLE,
				i_SIG => i_SIG,
				i_COEFF => i_COEFF,
				o_DFT => o_DFT,
				o_NEW_RESULT => o_NEW_RESULT
			 );
	
	
	   -- Clock process definitions
   i_clk_process :process
   begin
		i_CLK<= '0';
		wait for c_clk_period/2;
		i_CLK <= '1';
		wait for c_clk_period/2;
   end process;
	
	   -- Stimulus process
   stim_proc: process
	  variable L_IN : line;
	  variable CHAR : character;
	  variable DATA : std_logic_vector(7 downto 0);
	  file STIM_IN : text is in
						 "sine.dat";
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		i_ENABLE <= '1'; 
		i_COEFF <= to_signed(-2, CALC_WIDTH);
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
				i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(-1, INPUT_WIDTH);
		wait for signal_period/4;
		i_SIG <= to_signed(0, INPUT_WIDTH);
		wait for signal_period/4;
		-- File I/O signal gen
--		while not endfile(STIM_IN) loop
--			 readline(STIM_IN, L_IN);
--			 hread(L_IN, DATA);
--			 i_SIG <= signed(DATA);
--			 wait for signal_period;
--		end loop;
		
		wait;
		
   end process;
END;