--
--	Package File
--
--	Purpose: This package defines constants for AoA estimator

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package constants is

-- Declare constants

end constants;

package body constants is
 
end constants;
